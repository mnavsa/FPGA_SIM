library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity SEC is
port( 	CLK 			: in std_logic;
		PARITY_IN 		: in std_logic_vector(2 downto 0);
		CODEWORD_IN 	: in std_logic_vector(7 downto 0);
		CODEWORD_OUT 	: out std_logic_vector(7 downto 0);
		CORRECTED 		: out std_logic);
end SEC;

architecture RTL of SEC is
signal t_CORRECTED : std_logic := '0';
begin
	process(CLK,CODEWORD_IN)
	begin
		if PARITY_IN = "001" then 
			CODEWORD_OUT(0) <= NOT CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1'; 
		elsif PARITY_IN = "010" then 
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= NOT CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1';
		elsif PARITY_IN = "011" then 
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= NOT CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1';
		elsif PARITY_IN = "100" then 
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= NOT CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1';
		elsif PARITY_IN = "101" then 
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= NOT CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1';
		elsif PARITY_IN = "110" then 
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= NOT CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1';
		elsif PARITY_IN = "111" then 
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= NOT CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '1';
		else
			CODEWORD_OUT(0) <= CODEWORD_IN(0);
			CODEWORD_OUT(1) <= CODEWORD_IN(1);
			CODEWORD_OUT(2) <= CODEWORD_IN(2);
			CODEWORD_OUT(3) <= CODEWORD_IN(3);
			CODEWORD_OUT(4) <= CODEWORD_IN(4);
			CODEWORD_OUT(5) <= CODEWORD_IN(5);
			CODEWORD_OUT(6) <= CODEWORD_IN(6);
			CODEWORD_OUT(7) <= CODEWORD_IN(7);
			t_CORRECTED <= '0';
		end if;
	end process;
	CORRECTED <= t_CORRECTED;
end RTL;